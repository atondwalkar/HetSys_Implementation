module ast_data_cache_2w_v	(Resetn, MEM_address, MEM_in, WR, Clock, MEM_out, Done, RAM_addr_out, RAM_clk_out, RAM_inputdata_out, RAM_wen_out, RAM_outputdata_in, snoop_addr, snoop_wen, snoop_data);

//----------------------------------------------------------------------------
// 2-Way Set Associative Mapped Cache and Memory;
// The maximum memory capacity is 2^16 16-bit words.
// There are 2^5=32 words per block, and therefore 2^11 total blocks in MEM.
// The cache has 32 block locations.
// The address structure is: TAG=7-bit | Group=4-bit | Word=5-bit
// Two CAMs are used for each of the two ways.
// WR = 0 ==> READ; WR = 1 ==> WRITE.
//----------------------------------------------------------------------------

//----------------------------------------------------------------------------
// module parameters:
// ma_max = memory address width; md_max = memory data width;
// ca_max = cache address width; cam_addrs_max = cam address width;
// cam_arg_max = cam location/data width; cam_depth_max = total cam locations
// transfer count = 2^t_cnt = words per block
//----------------------------------------------------------------------------

//parameter ma_max=16, md_max=16, ca_max=10, t_cnt_max=5;
//parameter cam_addrs_max=4, cam_arg_max=7, cam_depth_max=16;

parameter ma_max=14, md_max=14, ca_max=7, t_cnt_max=4;
parameter cam_addrs_max=2, cam_arg_max=8, cam_depth_max=4;
parameter initfile = "blank.mif";

//----------------------------------------------------------------------------
// module input and output ports
//----------------------------------------------------------------------------
input [ma_max-1:0] MEM_address; // To speedup synthesis and simulation
input Resetn, WR, Clock;			// only 12K are being instantiated
input [md_max-1:0] MEM_in;
output [md_max-1:0] MEM_out;
output reg Done; // Means READ or WRITE ACCESS is complete, i.e. the output is 
	// valid during a READ, and done updating location during a WRITE
	
output [ma_max-1:0] RAM_addr_out;
output RAM_clk_out, RAM_wen_out;
output [md_max-1:0] RAM_inputdata_out;
input [md_max-1:0] RAM_outputdata_in;

input snoop_wen;
input [ma_max-1:0] snoop_addr;
input [md_max-1:0] snoop_data;
	
//----------------------------------------------------------------------------
// structural nets
//----------------------------------------------------------------------------
wire 	[cam_depth_max-1:0] mbits0, mbits1, grp;
wire	[md_max-1:0] MEMint_out, CACHE_out, CACHE_in;
wire	c0, c1, c2; // clock signals generated by the PLL
wire  	mem_clk, cache_clk;
wire	[cam_arg_max-1:0] dout0, dout1;
wire	[ma_max-1:0] MEMint_address; // internal memory address port
wire 	valid_snoop;
wire [ma_max-1:0] MEM_address_mux;

//----------------------------------------------------------------------------
// registered nets
//----------------------------------------------------------------------------
reg	[ma_max-1:0] MEMint_RDaddress, MEMint_WRaddress; // internal memory
reg	we0, we1, WRint, writeback;	// adress sources
reg	miss, wren, hit0, hit1;
reg [cam_depth_max-1:0] replace = {cam_depth_max{1'b0}};
reg	[ca_max-1:0] CACHE_address; // cache memory address	
reg	[cam_arg_max-1:0] din0, din1;
reg	[t_cnt_max:0] transfer_count;
reg	[cam_depth_max-1:0] cam0_init, cam1_init; // to mark the first upload
									// of a block of data to each cache block location
reg	[cam_depth_max-1:0] cam0_dirty_bit, cam1_dirty_bit; // to record if
reg 	[ma_max-1:0] MEM_snooped;
reg	snoop_status;
									// the block was ever written while in the cache 
//----------------------------------------------------------------------------
// grp_addrs_field is used to capture the value of the group address field
//----------------------------------------------------------------------------
integer	grp_addrs_field;
//----------------------------------------------------------------------------
// 7-bit Block Address | 4-bit Group Address | 5-bit Word Address
//----------------------------------------------------------------------------
// Structural part of the code = memory subsystem "data path"
//----------------------------------------------------------------------------
// The PLL unit/block generates three clock phases to sequence all events
//----------------------------------------------------------------------------
	ast_pll_3_v	my_pll 	(Clock, c0, c1, c2);
//----------------------------------------------------------------------------
// I'm using two separate CAM memories for the two-way TAG identification
//----------------------------------------------------------------------------
	//ast_CAM_v	my_cam0	(we0, 1'b1, din0, MEM_address_mux[ma_max-5:6], MEM_address_mux[5:4], dout0, mbits0);
	//ast_CAM_v	my_cam1	(we1, 1'b1, din1, MEM_address_mux[ma_max-5:6], MEM_address_mux[5:4], dout1, mbits1);
	
	assign valid_snoop = (snoop_wen && (&snoop_addr[13:8])); 
	
	assign MEM_address_mux = valid_snoop ? snoop_addr : MEM_address;
	
	ast_CAM_v	my_cam0	(we0, 1'b1, din0, MEM_address_mux[ma_max-1:6], MEM_address_mux[5:4], dout0, mbits0);
	ast_CAM_v	my_cam1	(we1, 1'b1, din1, MEM_address_mux[ma_max-1:6], MEM_address_mux[5:4], dout1, mbits1);
//----------------------------------------------------------------------------
// This is the actual MEM; an intitialized RAM; the same one that was used 
// before as a monolithic memory; notice that for a READ access this is driven
// by the c1 phase of the clock, while for a WRITE access by c2.
//----------------------------------------------------------------------------
	assign mem_clk = WRint ? c2 : c1;
	assign MEMint_address = writeback ? MEMint_WRaddress : MEMint_RDaddress;
	//astRISC521_ram1	my_ram	(MEMint_address[ma_max-5:0], mem_clk, CACHE_out, WRint, MEMint_out);
	//astRISC621_ram	#(.initfile(initfile)) my_ram	(MEMint_address[ma_max-1:0], mem_clk, CACHE_out, WRint, MEMint_out);
	assign RAM_addr_out = MEMint_address;
	assign RAM_clk_out = mem_clk;
	assign RAM_wen_out = WRint;
	assign RAM_inputdata_out = CACHE_out;
	assign MEMint_out = RAM_outputdata_in;
	//defparam prog_cache.my_ram.inifile = "file.mif";
//----------------------------------------------------------------------------
// This is the actual cache memory, implemented as a RAM; notice that for a 
// READ access this is driven by the c2 phase of the clock, while for a WRITE
// access by c1.
//----------------------------------------------------------------------------
	assign cache_clk = WRint ? c1 : c2;
	assign CACHE_in = valid_snoop ? snoop_data : (((hit0 || hit1) && WR) ? MEM_in : MEMint_out);
	//ast_cache_v			my_cache	(CACHE_address, cache_clk, CACHE_in, wren, CACHE_out);
	ast_cache_v			my_cache	(CACHE_address, cache_clk, CACHE_in, wren, CACHE_out);
	assign MEM_out = Done ? CACHE_out : {md_max{1'bz}};
//----------------------------------------------------------------------------
// This 4to16 decoder identifies the group being accessed
//----------------------------------------------------------------------------
	//ast_4to16_dec	my_dec	(MEM_address_mux[5:4], grp);
	ast_2to4_dec	my_dec	(MEM_address_mux[5:4], grp);
//----------------------------------------------------------------------------
// Behavioral part of the code = memory subsystem "control unit"
//----------------------------------------------------------------------------


always @ (posedge c0) begin
	if (Resetn == 0) begin
//----------------------------------------------------------------------------
// Memory subsystem initialization; after a reset the cache content is
//    random, and thus the miss signal is set to 1; this in turn will trigger
//    the transfer of the first block from MEM into the cache.
//----------------------------------------------------------------------------
		miss = 1'b1; transfer_count = {(t_cnt_max+1){1'b0}}; replace = 4'b0000;
		we0 = 0; we1 = 0; hit0 = 0; hit1 = 0; Done = 0; WRint = 0;
		cam0_init[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
		cam1_init[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
		cam0_dirty_bit[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
		cam1_dirty_bit[cam_depth_max-1:0] = {cam_depth_max{1'b0}};
		snoop_status = 0;
		end
	else begin 	
	grp_addrs_field = MEM_address_mux[5:4];
	
	
		if(valid_snoop)
		begin
			if(|(mbits0 & grp & cam0_init))
			begin
				miss = 1;
				snoop_status = 1;
				replace[grp_addrs_field] = 1'b0;
			end
			else if (|(mbits1 & grp & cam1_init))
			begin
				miss = 1;
				snoop_status = 1;
				replace[grp_addrs_field] = 1'b1;
			end
			else
				miss = 0;
		end
		else
		begin
	//----------------------------------------------------------------------------
	// The HIT if statements
	//----------------------------------------------------------------------------
	// miss == 0 means we execute these statements under the assumption that we
	//    have not yet discovered a miss.
	//----------------------------------------------------------------------------
			if (miss == 0) begin
				we0 = 0; we1 = 0; hit0 = 0; hit1 = 0; Done = 0; WRint = 0; wren = 0;
	//----------------------------------------------------------------------------
	// The condition logically ANDs each mbit with the coresponding group line;
	// Then, all are logically OR-ed using the OR reduction operator.
	//----------------------------------------------------------------------------
				if (|(mbits0 & grp & cam0_init)) begin
	//----------------------------------------------------------------------------
	// Concatenated group and word address fields.
	//----------------------------------------------------------------------------
					CACHE_address = {1'b0, MEM_address_mux[5:0]}; 
					if (WR == 1) 
					begin 
						cam0_dirty_bit[grp_addrs_field] = 1; 
						wren = 1; 
					end 
					else 
					begin 
						wren = 0; 
					end
					//if(snoop_wen && (&snoop_addr[13:8])) begin miss = 1; transfer_count = {(t_cnt_max+1){1'b0}}; end
					//else begin 
					hit0 = 1; Done = 1; 
	//----------------------------------------------------------------------------
	// Apply the replacing strategy: if this block was accessed now and a 
	//    replacement will be necessary next, replace the other block.
	//----------------------------------------------------------------------------
					replace[grp_addrs_field] = 1'b1;	end
				else if (|(mbits1 & grp & cam1_init)) begin
	//----------------------------------------------------------------------------
	// Concatenated group and word address fields.
	//----------------------------------------------------------------------------
					CACHE_address = {1'b1, MEM_address_mux[5:0]}; 
					if (WR == 1) 
					begin
						cam1_dirty_bit[grp_addrs_field] = 1; 
						wren = 1; 
					end 
					else 
					begin 
						wren =0; 
					end
					//if(snoop_wen && (&snoop_addr[13:8])) begin miss = 1; transfer_count = {(t_cnt_max+1){1'b0}}; end
					//else begin 
					hit1 = 1; Done = 1; 
	//----------------------------------------------------------------------------
	// Apply the replacing strategy: if this block was accessed now and a 
	//    replacement will be necessary next, replace the other block.
	//----------------------------------------------------------------------------
					replace[grp_addrs_field] = 1'b0;	end
	//----------------------------------------------------------------------------
	// A miss has been discovered, and thus the MISS statements are executed next
	//----------------------------------------------------------------------------
			else begin miss = 1'b1; //transfer_count = {(t_cnt_max+1){1'b0}}; 
				end
		end
	end
//----------------------------------------------------------------------------
// The WRITEBACK if statements
// are executed if the dirty bit of the block to be replaced has been set
//----------------------------------------------------------------------------
		writeback = (miss &  
				((~replace[grp_addrs_field] & cam0_dirty_bit[grp_addrs_field]) 
				| (replace[grp_addrs_field] & cam1_dirty_bit[grp_addrs_field])));
		if (writeback == 1)
			begin wren = 1'b0;  we0 = 0; we1 = 0; WRint = 1;
//----------------------------------------------------------------------------
// The CACHE_address is equal to the concatenation of the replace[i] bit, the 
//    group address field, and the word address; replace[i] is 0 or 1, and is
//    actually implementing a very simple replacement strategy: replace the 
//    block that was not used last of the two blocks in the cache.
//----------------------------------------------------------------------------
			CACHE_address = {replace[grp_addrs_field], MEM_address_mux[5:4], transfer_count[3:0]};
//----------------------------------------------------------------------------
// The MEMint_WRaddress is equal to the entire address generated by the CPU
//----------------------------------------------------------------------------
			if (replace[grp_addrs_field] == 0) 
			MEMint_WRaddress = {dout0, MEM_address_mux[5:4], transfer_count[3:0]};
			else MEMint_WRaddress = {dout1, MEM_address_mux[5:4], transfer_count[3:0]};		
//----------------------------------------------------------------------------
// The word address is incremented by 1 to point to the next word in the block
//----------------------------------------------------------------------------
			transfer_count = transfer_count + 1'b1; 
//----------------------------------------------------------------------------
// Check for the end of the block writeback and reset the dirty bit
//----------------------------------------------------------------------------
			if (transfer_count == 5'b10001) begin
				transfer_count = {(t_cnt_max+1){1'b0}}; // writeback = 1;
					if (replace[grp_addrs_field] == 0) 
							cam0_dirty_bit[grp_addrs_field] = 0;
					else	cam1_dirty_bit[grp_addrs_field] = 0; 
			end			
		end			
//----------------------------------------------------------------------------
// The MISS if statements - upload requested block in the cache
//----------------------------------------------------------------------------
		if (miss == 1 && writeback == 0) begin
//----------------------------------------------------------------------------
// The CACHE_address is equal to the concatenation of the replace[i] bit, the 
//    group address field, and the word address; replace[i] is 0 or 1, and is
//    actually implementing a very simple replacement strategy: replace the 
//    block that was not used last of the two blocks in the cache.
//----------------------------------------------------------------------------
			CACHE_address = {replace[grp_addrs_field], MEM_address_mux[5:4], transfer_count[3:0]};
//----------------------------------------------------------------------------
// The MEMint_RDaddress is equal to the entire address generated by the CPU
//----------------------------------------------------------------------------
			MEMint_RDaddress = {MEM_address_mux[ma_max-1:4], transfer_count[3:0]};
//----------------------------------------------------------------------------
// This wren enables the writing of the next word into the cache.
//----------------------------------------------------------------------------
			wren = 1'b1; WRint = 0;
//----------------------------------------------------------------------------
// The word address is incremented by 1 to point to the next word in the block
//----------------------------------------------------------------------------
			transfer_count = transfer_count + 1'b1; // end
//----------------------------------------------------------------------------
// At the end of a block transfer, update the CAMs
//----------------------------------------------------------------------------
		if(snoop_status == 1 && valid_snoop == 0)
		begin
			snoop_status = 0;
			transfer_count = 5'b10001;
		end

		if (transfer_count == 5'b10001) begin
			miss = 0; wren = 0; transfer_count = 5'b00000;
			if (replace[grp_addrs_field] == 0) begin
//----------------------------------------------------------------------------
// din0 OR din1 is the TAG of the new block, and their location in the cam  
//    is determined in the structural part above by the grp_addrs_field value.
//----------------------------------------------------------------------------
				din0 = MEM_address_mux[ma_max-1:6]; we0 = 1; 
				if (cam0_init[grp_addrs_field] == 0)  cam0_init[grp_addrs_field] =1;
				end // This block location has been initialized after reset
			else begin
				din1 = MEM_address_mux[ma_max-1:6]; we1 = 1;
				if (cam1_init[grp_addrs_field] == 0)  cam1_init[grp_addrs_field] =1;
				end // This block location has been initialized after reset
		end
	end
end
end
endmodule
